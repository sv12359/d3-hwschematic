module slice0(input [8-1:0] in, output out);
  assign out = in[3];
endmodule
